--------------------------------------------------------------------------------
-- Project     : ESS FPGA Framework
--------------------------------------------------------------------------------
-- File        : register_bank_config_pkg.vhdl
-- Authors     : Christian Amstutz
-- Created     : 2018-03-14
-- Last update : 2018-05-28
-- Platform    :
-- Standard    : VHDL'93
--------------------------------------------------------------------------------
-- Description :
-- Problems    :
--------------------------------------------------------------------------------
-- Copyright (c) 2018 European Spallation Source ERIC
--------------------------------------------------------------------------------
-- Revisions   :
--
-- 0.01 : 2018-05-28  Christian Amstutz
--        Created
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

package register_bank_config is

  constant ADDRESS_WIDTH         : integer   := 16;
  constant REGISTER_WIDTH        : integer   := 32;
  constant UNDEFINED_FIELD_VALUE : std_logic := '0';

  -- register_write_en_t
  type register_write_en_t is record
     Control              : std_logic;
     IrqFlag              : std_logic;
     IrqEnable            : std_logic;
     PulseIrqMap          : std_logic;
     SWEvent              : std_logic;
     DataBufCtrl          : std_logic;
     TXDataBufCtrl        : std_logic;
     TxSegBufCtrl         : std_logic;
     EvCntPresc           : std_logic;
     UsecDivider          : std_logic;
     ClockControl         : std_logic;
     GPIODir              : std_logic;
     GPIOIn               : std_logic;
     GPIOOut              : std_logic;
     DCTarget             : std_logic;
     SeqRamCtrl           : std_logic;
     Prescaler0           : std_logic;
     Prescaler1           : std_logic;
     Prescaler2           : std_logic;
     Prescaler3           : std_logic;
     Prescaler4           : std_logic;
     Prescaler5           : std_logic;
     Prescaler6           : std_logic;
     Prescaler7           : std_logic;
     PrescPhase0          : std_logic;
     PrescPhase1          : std_logic;
     PrescPhase2          : std_logic;
     PrescPhase3          : std_logic;
     PrescPhase4          : std_logic;
     PrescPhase5          : std_logic;
     PrescPhase6          : std_logic;
     PrescPhase7          : std_logic;
     PrescTrig0           : std_logic;
     PrescTrig1           : std_logic;
     PrescTrig2           : std_logic;
     PrescTrig3           : std_logic;
     PrescTrig4           : std_logic;
     PrescTrig5           : std_logic;
     PrescTrig6           : std_logic;
     PrescTrig7           : std_logic;
     DBusTrig0            : std_logic;
     DBusTrig1            : std_logic;
     DBusTrig2            : std_logic;
     DBusTrig3            : std_logic;
     DBusTrig4            : std_logic;
     DBusTrig5            : std_logic;
     DBusTrig6            : std_logic;
     DBusTrig7            : std_logic;
     Pulse0Ctrl           : std_logic;
     Pulse0Presc          : std_logic;
     Pulse0Delay          : std_logic;
     Pulse0Width          : std_logic;
     Pulse1Ctrl           : std_logic;
     Pulse1Presc          : std_logic;
     Pulse1Delay          : std_logic;
     Pulse1Width          : std_logic;
     Pulse2Ctrl           : std_logic;
     Pulse2Presc          : std_logic;
     Pulse2Delay          : std_logic;
     Pulse2Width          : std_logic;
     Pulse3Ctrl           : std_logic;
     Pulse3Presc          : std_logic;
     Pulse3Delay          : std_logic;
     Pulse3Width          : std_logic;
     Pulse4Ctrl           : std_logic;
     Pulse4Presc          : std_logic;
     Pulse4Delay          : std_logic;
     Pulse4Width          : std_logic;
     Pulse5Ctrl           : std_logic;
     Pulse5Presc          : std_logic;
     Pulse5Delay          : std_logic;
     Pulse5Width          : std_logic;
     Pulse6Ctrl           : std_logic;
     Pulse6Presc          : std_logic;
     Pulse6Delay          : std_logic;
     Pulse6Width          : std_logic;
     Pulse7Ctrl           : std_logic;
     Pulse7Presc          : std_logic;
     Pulse7Delay          : std_logic;
     Pulse7Width          : std_logic;
     Pulse8Ctrl           : std_logic;
     Pulse8Presc          : std_logic;
     Pulse8Delay          : std_logic;
     Pulse8Width          : std_logic;
     Pulse9Ctrl           : std_logic;
     Pulse9Presc          : std_logic;
     Pulse9Delay          : std_logic;
     Pulse9Width          : std_logic;
     Pulse10Ctrl          : std_logic;
     Pulse10Presc         : std_logic;
     Pulse10Delay         : std_logic;
     Pulse10Width         : std_logic;
     Pulse11Ctrl          : std_logic;
     Pulse11Presc         : std_logic;
     Pulse11Delay         : std_logic;
     Pulse11Width         : std_logic;
     Pulse12Ctrl          : std_logic;
     Pulse12Presc         : std_logic;
     Pulse12Delay         : std_logic;
     Pulse12Width         : std_logic;
     Pulse13Ctrl          : std_logic;
     Pulse13Presc         : std_logic;
     Pulse13Delay         : std_logic;
     Pulse13Width         : std_logic;
     Pulse14Ctrl          : std_logic;
     Pulse14Presc         : std_logic;
     Pulse14Delay         : std_logic;
     Pulse14Width         : std_logic;
     Pulse15Ctrl          : std_logic;
     Pulse15Presc         : std_logic;
     Pulse15Delay         : std_logic;
     Pulse15Width         : std_logic;
     Pulse16Ctrl          : std_logic;
     Pulse16Presc         : std_logic;
     Pulse16Delay         : std_logic;
     Pulse16Width         : std_logic;
     Pulse17Ctrl          : std_logic;
     Pulse17Presc         : std_logic;
     Pulse17Delay         : std_logic;
     Pulse17Width         : std_logic;
     Pulse18Ctrl          : std_logic;
     Pulse18Presc         : std_logic;
     Pulse18Delay         : std_logic;
     Pulse18Width         : std_logic;
     Pulse19Ctrl          : std_logic;
     Pulse19Presc         : std_logic;
     Pulse19Delay         : std_logic;
     Pulse19Width         : std_logic;
     Pulse20Ctrl          : std_logic;
     Pulse20Presc         : std_logic;
     Pulse20Delay         : std_logic;
     Pulse20Width         : std_logic;
     Pulse21Ctrl          : std_logic;
     Pulse21Presc         : std_logic;
     Pulse21Delay         : std_logic;
     Pulse21Width         : std_logic;
     Pulse22Ctrl          : std_logic;
     Pulse22Presc         : std_logic;
     Pulse22Delay         : std_logic;
     Pulse22Width         : std_logic;
     Pulse23Ctrl          : std_logic;
     Pulse23Presc         : std_logic;
     Pulse23Delay         : std_logic;
     Pulse23Width         : std_logic;
     Pulse24Ctrl          : std_logic;
     Pulse24Presc         : std_logic;
     Pulse24Delay         : std_logic;
     Pulse24Width         : std_logic;
     Pulse25Ctrl          : std_logic;
     Pulse25Presc         : std_logic;
     Pulse25Delay         : std_logic;
     Pulse25Width         : std_logic;
     Pulse26Ctrl          : std_logic;
     Pulse26Presc         : std_logic;
     Pulse26Delay         : std_logic;
     Pulse26Width         : std_logic;
     Pulse27Ctrl          : std_logic;
     Pulse27Presc         : std_logic;
     Pulse27Delay         : std_logic;
     Pulse27Width         : std_logic;
     Pulse28Ctrl          : std_logic;
     Pulse28Presc         : std_logic;
     Pulse28Delay         : std_logic;
     Pulse28Width         : std_logic;
     Pulse29Ctrl          : std_logic;
     Pulse29Presc         : std_logic;
     Pulse29Delay         : std_logic;
     Pulse29Width         : std_logic;
     Pulse30Ctrl          : std_logic;
     Pulse30Presc         : std_logic;
     Pulse30Delay         : std_logic;
     Pulse30Width         : std_logic;
     Pulse31Ctrl          : std_logic;
     Pulse31Presc         : std_logic;
     Pulse31Delay         : std_logic;
     Pulse31Width         : std_logic;
     ESSControl           : std_logic;
  end record;

  -- field_write_en_t
  type field_write_en_t is record
     Control              : std_logic;
     IrqFlag              : std_logic;
     IrqEnable            : std_logic;
     PulseIrqMap          : std_logic;
     SWEvent              : std_logic;
     DataBufCtrl          : std_logic;
     TXDataBufCtrl        : std_logic;
     TxSegBufCtrl         : std_logic;
     EvCntPresc           : std_logic;
     UsecDivider          : std_logic;
     ClockControl         : std_logic;
     GPIODir              : std_logic;
     GPIOIn               : std_logic;
     GPIOOut              : std_logic;
     DCTarget             : std_logic;
     SeqRamCtrl           : std_logic;
     Prescaler0           : std_logic;
     Prescaler1           : std_logic;
     Prescaler2           : std_logic;
     Prescaler3           : std_logic;
     Prescaler4           : std_logic;
     Prescaler5           : std_logic;
     Prescaler6           : std_logic;
     Prescaler7           : std_logic;
     PrescPhase0          : std_logic;
     PrescPhase1          : std_logic;
     PrescPhase2          : std_logic;
     PrescPhase3          : std_logic;
     PrescPhase4          : std_logic;
     PrescPhase5          : std_logic;
     PrescPhase6          : std_logic;
     PrescPhase7          : std_logic;
     PrescTrig0           : std_logic;
     PrescTrig1           : std_logic;
     PrescTrig2           : std_logic;
     PrescTrig3           : std_logic;
     PrescTrig4           : std_logic;
     PrescTrig5           : std_logic;
     PrescTrig6           : std_logic;
     PrescTrig7           : std_logic;
     DBusTrig0            : std_logic;
     DBusTrig1            : std_logic;
     DBusTrig2            : std_logic;
     DBusTrig3            : std_logic;
     DBusTrig4            : std_logic;
     DBusTrig5            : std_logic;
     DBusTrig6            : std_logic;
     DBusTrig7            : std_logic;
     Pulse0Ctrl           : std_logic;
     Pulse0Presc          : std_logic;
     Pulse0Delay          : std_logic;
     Pulse0Width          : std_logic;
     Pulse1Ctrl           : std_logic;
     Pulse1Presc          : std_logic;
     Pulse1Delay          : std_logic;
     Pulse1Width          : std_logic;
     Pulse2Ctrl           : std_logic;
     Pulse2Presc          : std_logic;
     Pulse2Delay          : std_logic;
     Pulse2Width          : std_logic;
     Pulse3Ctrl           : std_logic;
     Pulse3Presc          : std_logic;
     Pulse3Delay          : std_logic;
     Pulse3Width          : std_logic;
     Pulse4Ctrl           : std_logic;
     Pulse4Presc          : std_logic;
     Pulse4Delay          : std_logic;
     Pulse4Width          : std_logic;
     Pulse5Ctrl           : std_logic;
     Pulse5Presc          : std_logic;
     Pulse5Delay          : std_logic;
     Pulse5Width          : std_logic;
     Pulse6Ctrl           : std_logic;
     Pulse6Presc          : std_logic;
     Pulse6Delay          : std_logic;
     Pulse6Width          : std_logic;
     Pulse7Ctrl           : std_logic;
     Pulse7Presc          : std_logic;
     Pulse7Delay          : std_logic;
     Pulse7Width          : std_logic;
     Pulse8Ctrl           : std_logic;
     Pulse8Presc          : std_logic;
     Pulse8Delay          : std_logic;
     Pulse8Width          : std_logic;
     Pulse9Ctrl           : std_logic;
     Pulse9Presc          : std_logic;
     Pulse9Delay          : std_logic;
     Pulse9Width          : std_logic;
     Pulse10Ctrl          : std_logic;
     Pulse10Presc         : std_logic;
     Pulse10Delay         : std_logic;
     Pulse10Width         : std_logic;
     Pulse11Ctrl          : std_logic;
     Pulse11Presc         : std_logic;
     Pulse11Delay         : std_logic;
     Pulse11Width         : std_logic;
     Pulse12Ctrl          : std_logic;
     Pulse12Presc         : std_logic;
     Pulse12Delay         : std_logic;
     Pulse12Width         : std_logic;
     Pulse13Ctrl          : std_logic;
     Pulse13Presc         : std_logic;
     Pulse13Delay         : std_logic;
     Pulse13Width         : std_logic;
     Pulse14Ctrl          : std_logic;
     Pulse14Presc         : std_logic;
     Pulse14Delay         : std_logic;
     Pulse14Width         : std_logic;
     Pulse15Ctrl          : std_logic;
     Pulse15Presc         : std_logic;
     Pulse15Delay         : std_logic;
     Pulse15Width         : std_logic;
     Pulse16Ctrl          : std_logic;
     Pulse16Presc         : std_logic;
     Pulse16Delay         : std_logic;
     Pulse16Width         : std_logic;
     Pulse17Ctrl          : std_logic;
     Pulse17Presc         : std_logic;
     Pulse17Delay         : std_logic;
     Pulse17Width         : std_logic;
     Pulse18Ctrl          : std_logic;
     Pulse18Presc         : std_logic;
     Pulse18Delay         : std_logic;
     Pulse18Width         : std_logic;
     Pulse19Ctrl          : std_logic;
     Pulse19Presc         : std_logic;
     Pulse19Delay         : std_logic;
     Pulse19Width         : std_logic;
     Pulse20Ctrl          : std_logic;
     Pulse20Presc         : std_logic;
     Pulse20Delay         : std_logic;
     Pulse20Width         : std_logic;
     Pulse21Ctrl          : std_logic;
     Pulse21Presc         : std_logic;
     Pulse21Delay         : std_logic;
     Pulse21Width         : std_logic;
     Pulse22Ctrl          : std_logic;
     Pulse22Presc         : std_logic;
     Pulse22Delay         : std_logic;
     Pulse22Width         : std_logic;
     Pulse23Ctrl          : std_logic;
     Pulse23Presc         : std_logic;
     Pulse23Delay         : std_logic;
     Pulse23Width         : std_logic;
     Pulse24Ctrl          : std_logic;
     Pulse24Presc         : std_logic;
     Pulse24Delay         : std_logic;
     Pulse24Width         : std_logic;
     Pulse25Ctrl          : std_logic;
     Pulse25Presc         : std_logic;
     Pulse25Delay         : std_logic;
     Pulse25Width         : std_logic;
     Pulse26Ctrl          : std_logic;
     Pulse26Presc         : std_logic;
     Pulse26Delay         : std_logic;
     Pulse26Width         : std_logic;
     Pulse27Ctrl          : std_logic;
     Pulse27Presc         : std_logic;
     Pulse27Delay         : std_logic;
     Pulse27Width         : std_logic;
     Pulse28Ctrl          : std_logic;
     Pulse28Presc         : std_logic;
     Pulse28Delay         : std_logic;
     Pulse28Width         : std_logic;
     Pulse29Ctrl          : std_logic;
     Pulse29Presc         : std_logic;
     Pulse29Delay         : std_logic;
     Pulse29Width         : std_logic;
     Pulse30Ctrl          : std_logic;
     Pulse30Presc         : std_logic;
     Pulse30Delay         : std_logic;
     Pulse30Width         : std_logic;
     Pulse31Ctrl          : std_logic;
     Pulse31Presc         : std_logic;
     Pulse31Delay         : std_logic;
     Pulse31Width         : std_logic;
     ESSControl           : std_logic;
  end record;

  -- field_data_t
  type field_data_t is record
     Status               : std_logic_vector(31 downto 0);
     Control              : std_logic_vector(31 downto 0);
     IrqFlag              : std_logic_vector(31 downto 0);
     IrqEnable            : std_logic_vector(31 downto 0);
     PulseIrqMap          : std_logic_vector(31 downto 0);
     SWEvent              : std_logic_vector(31 downto 0);
     DataBufCtrl          : std_logic_vector(31 downto 0);
     TXDataBufCtrl        : std_logic_vector(31 downto 0);
     TxSegBufCtrl         : std_logic_vector(31 downto 0);
     FWVersion            : std_logic_vector(31 downto 0);
     EvCntPresc           : std_logic_vector(31 downto 0);
     UsecDivider          : std_logic_vector(31 downto 0);
     ClockControl         : std_logic_vector(31 downto 0);
     SecSR                : std_logic_vector(31 downto 0);
     SecCounter           : std_logic_vector(31 downto 0);
     EventCounter         : std_logic_vector(31 downto 0);
     SecLatch             : std_logic_vector(31 downto 0);
     EvCntLatch           : std_logic_vector(31 downto 0);
     EvFIFOSec            : std_logic_vector(31 downto 0);
     EvFIFOEvCnt          : std_logic_vector(31 downto 0);
     EvFIFOCode           : std_logic_vector(31 downto 0);
     LogStatus            : std_logic_vector(31 downto 0);
     GPIODir              : std_logic_vector(31 downto 0);
     GPIOIn               : std_logic_vector(31 downto 0);
     GPIOOut              : std_logic_vector(31 downto 0);
     DCTarget             : std_logic_vector(31 downto 0);
     DCRxValue            : std_logic_vector(31 downto 0);
     DCIntValue           : std_logic_vector(31 downto 0);
     DCStatus             : std_logic_vector(31 downto 0);
     TopologyID           : std_logic_vector(31 downto 0);
     SeqRamCtrl           : std_logic_vector(31 downto 0);
     Prescaler0           : std_logic_vector(31 downto 0);
     Prescaler1           : std_logic_vector(31 downto 0);
     Prescaler2           : std_logic_vector(31 downto 0);
     Prescaler3           : std_logic_vector(31 downto 0);
     Prescaler4           : std_logic_vector(31 downto 0);
     Prescaler5           : std_logic_vector(31 downto 0);
     Prescaler6           : std_logic_vector(31 downto 0);
     Prescaler7           : std_logic_vector(31 downto 0);
     PrescPhase0          : std_logic_vector(31 downto 0);
     PrescPhase1          : std_logic_vector(31 downto 0);
     PrescPhase2          : std_logic_vector(31 downto 0);
     PrescPhase3          : std_logic_vector(31 downto 0);
     PrescPhase4          : std_logic_vector(31 downto 0);
     PrescPhase5          : std_logic_vector(31 downto 0);
     PrescPhase6          : std_logic_vector(31 downto 0);
     PrescPhase7          : std_logic_vector(31 downto 0);
     PrescTrig0           : std_logic_vector(31 downto 0);
     PrescTrig1           : std_logic_vector(31 downto 0);
     PrescTrig2           : std_logic_vector(31 downto 0);
     PrescTrig3           : std_logic_vector(31 downto 0);
     PrescTrig4           : std_logic_vector(31 downto 0);
     PrescTrig5           : std_logic_vector(31 downto 0);
     PrescTrig6           : std_logic_vector(31 downto 0);
     PrescTrig7           : std_logic_vector(31 downto 0);
     DBusTrig0            : std_logic_vector(31 downto 0);
     DBusTrig1            : std_logic_vector(31 downto 0);
     DBusTrig2            : std_logic_vector(31 downto 0);
     DBusTrig3            : std_logic_vector(31 downto 0);
     DBusTrig4            : std_logic_vector(31 downto 0);
     DBusTrig5            : std_logic_vector(31 downto 0);
     DBusTrig6            : std_logic_vector(31 downto 0);
     DBusTrig7            : std_logic_vector(31 downto 0);
     Pulse0Ctrl           : std_logic_vector(31 downto 0);
     Pulse0Presc          : std_logic_vector(31 downto 0);
     Pulse0Delay          : std_logic_vector(31 downto 0);
     Pulse0Width          : std_logic_vector(31 downto 0);
     Pulse1Ctrl           : std_logic_vector(31 downto 0);
     Pulse1Presc          : std_logic_vector(31 downto 0);
     Pulse1Delay          : std_logic_vector(31 downto 0);
     Pulse1Width          : std_logic_vector(31 downto 0);
     Pulse2Ctrl           : std_logic_vector(31 downto 0);
     Pulse2Presc          : std_logic_vector(31 downto 0);
     Pulse2Delay          : std_logic_vector(31 downto 0);
     Pulse2Width          : std_logic_vector(31 downto 0);
     Pulse3Ctrl           : std_logic_vector(31 downto 0);
     Pulse3Presc          : std_logic_vector(31 downto 0);
     Pulse3Delay          : std_logic_vector(31 downto 0);
     Pulse3Width          : std_logic_vector(31 downto 0);
     Pulse4Ctrl           : std_logic_vector(31 downto 0);
     Pulse4Presc          : std_logic_vector(31 downto 0);
     Pulse4Delay          : std_logic_vector(31 downto 0);
     Pulse4Width          : std_logic_vector(31 downto 0);
     Pulse5Ctrl           : std_logic_vector(31 downto 0);
     Pulse5Presc          : std_logic_vector(31 downto 0);
     Pulse5Delay          : std_logic_vector(31 downto 0);
     Pulse5Width          : std_logic_vector(31 downto 0);
     Pulse6Ctrl           : std_logic_vector(31 downto 0);
     Pulse6Presc          : std_logic_vector(31 downto 0);
     Pulse6Delay          : std_logic_vector(31 downto 0);
     Pulse6Width          : std_logic_vector(31 downto 0);
     Pulse7Ctrl           : std_logic_vector(31 downto 0);
     Pulse7Presc          : std_logic_vector(31 downto 0);
     Pulse7Delay          : std_logic_vector(31 downto 0);
     Pulse7Width          : std_logic_vector(31 downto 0);
     Pulse8Ctrl           : std_logic_vector(31 downto 0);
     Pulse8Presc          : std_logic_vector(31 downto 0);
     Pulse8Delay          : std_logic_vector(31 downto 0);
     Pulse8Width          : std_logic_vector(31 downto 0);
     Pulse9Ctrl           : std_logic_vector(31 downto 0);
     Pulse9Presc          : std_logic_vector(31 downto 0);
     Pulse9Delay          : std_logic_vector(31 downto 0);
     Pulse9Width          : std_logic_vector(31 downto 0);
     Pulse10Ctrl          : std_logic_vector(31 downto 0);
     Pulse10Presc         : std_logic_vector(31 downto 0);
     Pulse10Delay         : std_logic_vector(31 downto 0);
     Pulse10Width         : std_logic_vector(31 downto 0);
     Pulse11Ctrl          : std_logic_vector(31 downto 0);
     Pulse11Presc         : std_logic_vector(31 downto 0);
     Pulse11Delay         : std_logic_vector(31 downto 0);
     Pulse11Width         : std_logic_vector(31 downto 0);
     Pulse12Ctrl          : std_logic_vector(31 downto 0);
     Pulse12Presc         : std_logic_vector(31 downto 0);
     Pulse12Delay         : std_logic_vector(31 downto 0);
     Pulse12Width         : std_logic_vector(31 downto 0);
     Pulse13Ctrl          : std_logic_vector(31 downto 0);
     Pulse13Presc         : std_logic_vector(31 downto 0);
     Pulse13Delay         : std_logic_vector(31 downto 0);
     Pulse13Width         : std_logic_vector(31 downto 0);
     Pulse14Ctrl          : std_logic_vector(31 downto 0);
     Pulse14Presc         : std_logic_vector(31 downto 0);
     Pulse14Delay         : std_logic_vector(31 downto 0);
     Pulse14Width         : std_logic_vector(31 downto 0);
     Pulse15Ctrl          : std_logic_vector(31 downto 0);
     Pulse15Presc         : std_logic_vector(31 downto 0);
     Pulse15Delay         : std_logic_vector(31 downto 0);
     Pulse15Width         : std_logic_vector(31 downto 0);
     Pulse16Ctrl          : std_logic_vector(31 downto 0);
     Pulse16Presc         : std_logic_vector(31 downto 0);
     Pulse16Delay         : std_logic_vector(31 downto 0);
     Pulse16Width         : std_logic_vector(31 downto 0);
     Pulse17Ctrl          : std_logic_vector(31 downto 0);
     Pulse17Presc         : std_logic_vector(31 downto 0);
     Pulse17Delay         : std_logic_vector(31 downto 0);
     Pulse17Width         : std_logic_vector(31 downto 0);
     Pulse18Ctrl          : std_logic_vector(31 downto 0);
     Pulse18Presc         : std_logic_vector(31 downto 0);
     Pulse18Delay         : std_logic_vector(31 downto 0);
     Pulse18Width         : std_logic_vector(31 downto 0);
     Pulse19Ctrl          : std_logic_vector(31 downto 0);
     Pulse19Presc         : std_logic_vector(31 downto 0);
     Pulse19Delay         : std_logic_vector(31 downto 0);
     Pulse19Width         : std_logic_vector(31 downto 0);
     Pulse20Ctrl          : std_logic_vector(31 downto 0);
     Pulse20Presc         : std_logic_vector(31 downto 0);
     Pulse20Delay         : std_logic_vector(31 downto 0);
     Pulse20Width         : std_logic_vector(31 downto 0);
     Pulse21Ctrl          : std_logic_vector(31 downto 0);
     Pulse21Presc         : std_logic_vector(31 downto 0);
     Pulse21Delay         : std_logic_vector(31 downto 0);
     Pulse21Width         : std_logic_vector(31 downto 0);
     Pulse22Ctrl          : std_logic_vector(31 downto 0);
     Pulse22Presc         : std_logic_vector(31 downto 0);
     Pulse22Delay         : std_logic_vector(31 downto 0);
     Pulse22Width         : std_logic_vector(31 downto 0);
     Pulse23Ctrl          : std_logic_vector(31 downto 0);
     Pulse23Presc         : std_logic_vector(31 downto 0);
     Pulse23Delay         : std_logic_vector(31 downto 0);
     Pulse23Width         : std_logic_vector(31 downto 0);
     Pulse24Ctrl          : std_logic_vector(31 downto 0);
     Pulse24Presc         : std_logic_vector(31 downto 0);
     Pulse24Delay         : std_logic_vector(31 downto 0);
     Pulse24Width         : std_logic_vector(31 downto 0);
     Pulse25Ctrl          : std_logic_vector(31 downto 0);
     Pulse25Presc         : std_logic_vector(31 downto 0);
     Pulse25Delay         : std_logic_vector(31 downto 0);
     Pulse25Width         : std_logic_vector(31 downto 0);
     Pulse26Ctrl          : std_logic_vector(31 downto 0);
     Pulse26Presc         : std_logic_vector(31 downto 0);
     Pulse26Delay         : std_logic_vector(31 downto 0);
     Pulse26Width         : std_logic_vector(31 downto 0);
     Pulse27Ctrl          : std_logic_vector(31 downto 0);
     Pulse27Presc         : std_logic_vector(31 downto 0);
     Pulse27Delay         : std_logic_vector(31 downto 0);
     Pulse27Width         : std_logic_vector(31 downto 0);
     Pulse28Ctrl          : std_logic_vector(31 downto 0);
     Pulse28Presc         : std_logic_vector(31 downto 0);
     Pulse28Delay         : std_logic_vector(31 downto 0);
     Pulse28Width         : std_logic_vector(31 downto 0);
     Pulse29Ctrl          : std_logic_vector(31 downto 0);
     Pulse29Presc         : std_logic_vector(31 downto 0);
     Pulse29Delay         : std_logic_vector(31 downto 0);
     Pulse29Width         : std_logic_vector(31 downto 0);
     Pulse30Ctrl          : std_logic_vector(31 downto 0);
     Pulse30Presc         : std_logic_vector(31 downto 0);
     Pulse30Delay         : std_logic_vector(31 downto 0);
     Pulse30Width         : std_logic_vector(31 downto 0);
     Pulse31Ctrl          : std_logic_vector(31 downto 0);
     Pulse31Presc         : std_logic_vector(31 downto 0);
     Pulse31Delay         : std_logic_vector(31 downto 0);
     Pulse31Width         : std_logic_vector(31 downto 0);
     ESSStatus            : std_logic_vector(31 downto 0);
     ESSControl           : std_logic_vector(31 downto 0);
     ESSExtSecCounter     : std_logic_vector(31 downto 0);
     ESSExtEventCounter   : std_logic_vector(31 downto 0);
  end record;

  -- register_bus_read_t
  type register_bus_read_t is record
     Status               : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Control              : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     IrqFlag              : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     IrqEnable            : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     PulseIrqMap          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     SWEvent              : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     DataBufCtrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     TXDataBufCtrl        : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     TxSegBufCtrl         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     FWVersion            : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     EvCntPresc           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     UsecDivider          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     ClockControl         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     SecSR                : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     SecCounter           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     EventCounter         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     SecLatch             : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     EvCntLatch           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     EvFIFOSec            : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     EvFIFOEvCnt          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     EvFIFOCode           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     LogStatus            : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     GPIODir              : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     GPIOIn               : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     GPIOOut              : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     DCTarget             : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     DCRxValue            : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     DCIntValue           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     DCStatus             : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     TopologyID           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     SeqRamCtrl           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Prescaler0           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Prescaler1           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Prescaler2           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Prescaler3           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Prescaler4           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Prescaler5           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Prescaler6           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Prescaler7           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     PrescPhase0          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     PrescPhase1          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     PrescPhase2          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     PrescPhase3          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     PrescPhase4          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     PrescPhase5          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     PrescPhase6          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     PrescPhase7          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     PrescTrig0           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     PrescTrig1           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     PrescTrig2           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     PrescTrig3           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     PrescTrig4           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     PrescTrig5           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     PrescTrig6           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     PrescTrig7           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     DBusTrig0            : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     DBusTrig1            : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     DBusTrig2            : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     DBusTrig3            : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     DBusTrig4            : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     DBusTrig5            : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     DBusTrig6            : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     DBusTrig7            : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse0Ctrl           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse0Presc          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse0Delay          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse0Width          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse1Ctrl           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse1Presc          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse1Delay          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse1Width          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse2Ctrl           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse2Presc          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse2Delay          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse2Width          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse3Ctrl           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse3Presc          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse3Delay          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse3Width          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse4Ctrl           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse4Presc          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse4Delay          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse4Width          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse5Ctrl           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse5Presc          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse5Delay          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse5Width          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse6Ctrl           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse6Presc          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse6Delay          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse6Width          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse7Ctrl           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse7Presc          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse7Delay          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse7Width          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse8Ctrl           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse8Presc          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse8Delay          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse8Width          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse9Ctrl           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse9Presc          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse9Delay          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse9Width          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse10Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse10Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse10Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse10Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse11Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse11Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse11Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse11Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse12Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse12Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse12Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse12Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse13Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse13Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse13Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse13Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse14Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse14Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse14Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse14Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse15Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse15Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse15Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse15Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse16Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse16Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse16Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse16Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse17Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse17Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse17Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse17Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse18Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse18Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse18Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse18Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse19Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse19Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse19Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse19Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse20Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse20Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse20Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse20Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse21Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse21Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse21Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse21Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse22Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse22Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse22Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse22Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse23Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse23Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse23Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse23Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse24Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse24Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse24Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse24Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse25Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse25Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse25Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse25Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse26Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse26Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse26Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse26Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse27Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse27Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse27Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse27Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse28Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse28Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse28Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse28Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse29Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse29Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse29Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse29Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse30Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse30Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse30Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse30Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse31Ctrl          : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse31Presc         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse31Delay         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     Pulse31Width         : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     ESSStatus            : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     ESSControl           : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     ESSExtSecCounter     : std_logic_vector(REGISTER_WIDTH-1 downto 0);
     ESSExtEventCounter   : std_logic_vector(REGISTER_WIDTH-1 downto 0);
  end record;

  -- logic_read_data_t
  type logic_read_data_t is record
     Control              : std_logic_vector(31 downto 0);
     IrqFlag              : std_logic_vector(31 downto 0);
     IrqEnable            : std_logic_vector(31 downto 0);
     PulseIrqMap          : std_logic_vector(31 downto 0);
     SWEvent              : std_logic_vector(31 downto 0);
     DataBufCtrl          : std_logic_vector(31 downto 0);
     TXDataBufCtrl        : std_logic_vector(31 downto 0);
     TxSegBufCtrl         : std_logic_vector(31 downto 0);
     EvCntPresc           : std_logic_vector(31 downto 0);
     UsecDivider          : std_logic_vector(31 downto 0);
     ClockControl         : std_logic_vector(31 downto 0);
     GPIODir              : std_logic_vector(31 downto 0);
     GPIOIn               : std_logic_vector(31 downto 0);
     GPIOOut              : std_logic_vector(31 downto 0);
     DCTarget             : std_logic_vector(31 downto 0);
     SeqRamCtrl           : std_logic_vector(31 downto 0);
     Prescaler0           : std_logic_vector(31 downto 0);
     Prescaler1           : std_logic_vector(31 downto 0);
     Prescaler2           : std_logic_vector(31 downto 0);
     Prescaler3           : std_logic_vector(31 downto 0);
     Prescaler4           : std_logic_vector(31 downto 0);
     Prescaler5           : std_logic_vector(31 downto 0);
     Prescaler6           : std_logic_vector(31 downto 0);
     Prescaler7           : std_logic_vector(31 downto 0);
     PrescPhase0          : std_logic_vector(31 downto 0);
     PrescPhase1          : std_logic_vector(31 downto 0);
     PrescPhase2          : std_logic_vector(31 downto 0);
     PrescPhase3          : std_logic_vector(31 downto 0);
     PrescPhase4          : std_logic_vector(31 downto 0);
     PrescPhase5          : std_logic_vector(31 downto 0);
     PrescPhase6          : std_logic_vector(31 downto 0);
     PrescPhase7          : std_logic_vector(31 downto 0);
     PrescTrig0           : std_logic_vector(31 downto 0);
     PrescTrig1           : std_logic_vector(31 downto 0);
     PrescTrig2           : std_logic_vector(31 downto 0);
     PrescTrig3           : std_logic_vector(31 downto 0);
     PrescTrig4           : std_logic_vector(31 downto 0);
     PrescTrig5           : std_logic_vector(31 downto 0);
     PrescTrig6           : std_logic_vector(31 downto 0);
     PrescTrig7           : std_logic_vector(31 downto 0);
     DBusTrig0            : std_logic_vector(31 downto 0);
     DBusTrig1            : std_logic_vector(31 downto 0);
     DBusTrig2            : std_logic_vector(31 downto 0);
     DBusTrig3            : std_logic_vector(31 downto 0);
     DBusTrig4            : std_logic_vector(31 downto 0);
     DBusTrig5            : std_logic_vector(31 downto 0);
     DBusTrig6            : std_logic_vector(31 downto 0);
     DBusTrig7            : std_logic_vector(31 downto 0);
     Pulse0Ctrl           : std_logic_vector(31 downto 0);
     Pulse0Presc          : std_logic_vector(31 downto 0);
     Pulse0Delay          : std_logic_vector(31 downto 0);
     Pulse0Width          : std_logic_vector(31 downto 0);
     Pulse1Ctrl           : std_logic_vector(31 downto 0);
     Pulse1Presc          : std_logic_vector(31 downto 0);
     Pulse1Delay          : std_logic_vector(31 downto 0);
     Pulse1Width          : std_logic_vector(31 downto 0);
     Pulse2Ctrl           : std_logic_vector(31 downto 0);
     Pulse2Presc          : std_logic_vector(31 downto 0);
     Pulse2Delay          : std_logic_vector(31 downto 0);
     Pulse2Width          : std_logic_vector(31 downto 0);
     Pulse3Ctrl           : std_logic_vector(31 downto 0);
     Pulse3Presc          : std_logic_vector(31 downto 0);
     Pulse3Delay          : std_logic_vector(31 downto 0);
     Pulse3Width          : std_logic_vector(31 downto 0);
     Pulse4Ctrl           : std_logic_vector(31 downto 0);
     Pulse4Presc          : std_logic_vector(31 downto 0);
     Pulse4Delay          : std_logic_vector(31 downto 0);
     Pulse4Width          : std_logic_vector(31 downto 0);
     Pulse5Ctrl           : std_logic_vector(31 downto 0);
     Pulse5Presc          : std_logic_vector(31 downto 0);
     Pulse5Delay          : std_logic_vector(31 downto 0);
     Pulse5Width          : std_logic_vector(31 downto 0);
     Pulse6Ctrl           : std_logic_vector(31 downto 0);
     Pulse6Presc          : std_logic_vector(31 downto 0);
     Pulse6Delay          : std_logic_vector(31 downto 0);
     Pulse6Width          : std_logic_vector(31 downto 0);
     Pulse7Ctrl           : std_logic_vector(31 downto 0);
     Pulse7Presc          : std_logic_vector(31 downto 0);
     Pulse7Delay          : std_logic_vector(31 downto 0);
     Pulse7Width          : std_logic_vector(31 downto 0);
     Pulse8Ctrl           : std_logic_vector(31 downto 0);
     Pulse8Presc          : std_logic_vector(31 downto 0);
     Pulse8Delay          : std_logic_vector(31 downto 0);
     Pulse8Width          : std_logic_vector(31 downto 0);
     Pulse9Ctrl           : std_logic_vector(31 downto 0);
     Pulse9Presc          : std_logic_vector(31 downto 0);
     Pulse9Delay          : std_logic_vector(31 downto 0);
     Pulse9Width          : std_logic_vector(31 downto 0);
     Pulse10Ctrl          : std_logic_vector(31 downto 0);
     Pulse10Presc         : std_logic_vector(31 downto 0);
     Pulse10Delay         : std_logic_vector(31 downto 0);
     Pulse10Width         : std_logic_vector(31 downto 0);
     Pulse11Ctrl          : std_logic_vector(31 downto 0);
     Pulse11Presc         : std_logic_vector(31 downto 0);
     Pulse11Delay         : std_logic_vector(31 downto 0);
     Pulse11Width         : std_logic_vector(31 downto 0);
     Pulse12Ctrl          : std_logic_vector(31 downto 0);
     Pulse12Presc         : std_logic_vector(31 downto 0);
     Pulse12Delay         : std_logic_vector(31 downto 0);
     Pulse12Width         : std_logic_vector(31 downto 0);
     Pulse13Ctrl          : std_logic_vector(31 downto 0);
     Pulse13Presc         : std_logic_vector(31 downto 0);
     Pulse13Delay         : std_logic_vector(31 downto 0);
     Pulse13Width         : std_logic_vector(31 downto 0);
     Pulse14Ctrl          : std_logic_vector(31 downto 0);
     Pulse14Presc         : std_logic_vector(31 downto 0);
     Pulse14Delay         : std_logic_vector(31 downto 0);
     Pulse14Width         : std_logic_vector(31 downto 0);
     Pulse15Ctrl          : std_logic_vector(31 downto 0);
     Pulse15Presc         : std_logic_vector(31 downto 0);
     Pulse15Delay         : std_logic_vector(31 downto 0);
     Pulse15Width         : std_logic_vector(31 downto 0);
     Pulse16Ctrl          : std_logic_vector(31 downto 0);
     Pulse16Presc         : std_logic_vector(31 downto 0);
     Pulse16Delay         : std_logic_vector(31 downto 0);
     Pulse16Width         : std_logic_vector(31 downto 0);
     Pulse17Ctrl          : std_logic_vector(31 downto 0);
     Pulse17Presc         : std_logic_vector(31 downto 0);
     Pulse17Delay         : std_logic_vector(31 downto 0);
     Pulse17Width         : std_logic_vector(31 downto 0);
     Pulse18Ctrl          : std_logic_vector(31 downto 0);
     Pulse18Presc         : std_logic_vector(31 downto 0);
     Pulse18Delay         : std_logic_vector(31 downto 0);
     Pulse18Width         : std_logic_vector(31 downto 0);
     Pulse19Ctrl          : std_logic_vector(31 downto 0);
     Pulse19Presc         : std_logic_vector(31 downto 0);
     Pulse19Delay         : std_logic_vector(31 downto 0);
     Pulse19Width         : std_logic_vector(31 downto 0);
     Pulse20Ctrl          : std_logic_vector(31 downto 0);
     Pulse20Presc         : std_logic_vector(31 downto 0);
     Pulse20Delay         : std_logic_vector(31 downto 0);
     Pulse20Width         : std_logic_vector(31 downto 0);
     Pulse21Ctrl          : std_logic_vector(31 downto 0);
     Pulse21Presc         : std_logic_vector(31 downto 0);
     Pulse21Delay         : std_logic_vector(31 downto 0);
     Pulse21Width         : std_logic_vector(31 downto 0);
     Pulse22Ctrl          : std_logic_vector(31 downto 0);
     Pulse22Presc         : std_logic_vector(31 downto 0);
     Pulse22Delay         : std_logic_vector(31 downto 0);
     Pulse22Width         : std_logic_vector(31 downto 0);
     Pulse23Ctrl          : std_logic_vector(31 downto 0);
     Pulse23Presc         : std_logic_vector(31 downto 0);
     Pulse23Delay         : std_logic_vector(31 downto 0);
     Pulse23Width         : std_logic_vector(31 downto 0);
     Pulse24Ctrl          : std_logic_vector(31 downto 0);
     Pulse24Presc         : std_logic_vector(31 downto 0);
     Pulse24Delay         : std_logic_vector(31 downto 0);
     Pulse24Width         : std_logic_vector(31 downto 0);
     Pulse25Ctrl          : std_logic_vector(31 downto 0);
     Pulse25Presc         : std_logic_vector(31 downto 0);
     Pulse25Delay         : std_logic_vector(31 downto 0);
     Pulse25Width         : std_logic_vector(31 downto 0);
     Pulse26Ctrl          : std_logic_vector(31 downto 0);
     Pulse26Presc         : std_logic_vector(31 downto 0);
     Pulse26Delay         : std_logic_vector(31 downto 0);
     Pulse26Width         : std_logic_vector(31 downto 0);
     Pulse27Ctrl          : std_logic_vector(31 downto 0);
     Pulse27Presc         : std_logic_vector(31 downto 0);
     Pulse27Delay         : std_logic_vector(31 downto 0);
     Pulse27Width         : std_logic_vector(31 downto 0);
     Pulse28Ctrl          : std_logic_vector(31 downto 0);
     Pulse28Presc         : std_logic_vector(31 downto 0);
     Pulse28Delay         : std_logic_vector(31 downto 0);
     Pulse28Width         : std_logic_vector(31 downto 0);
     Pulse29Ctrl          : std_logic_vector(31 downto 0);
     Pulse29Presc         : std_logic_vector(31 downto 0);
     Pulse29Delay         : std_logic_vector(31 downto 0);
     Pulse29Width         : std_logic_vector(31 downto 0);
     Pulse30Ctrl          : std_logic_vector(31 downto 0);
     Pulse30Presc         : std_logic_vector(31 downto 0);
     Pulse30Delay         : std_logic_vector(31 downto 0);
     Pulse30Width         : std_logic_vector(31 downto 0);
     Pulse31Ctrl          : std_logic_vector(31 downto 0);
     Pulse31Presc         : std_logic_vector(31 downto 0);
     Pulse31Delay         : std_logic_vector(31 downto 0);
     Pulse31Width         : std_logic_vector(31 downto 0);
     ESSControl           : std_logic_vector(31 downto 0);
  end record;

  -- logic_return_t
  type logic_return_t is record
     Status               : std_logic_vector(31 downto 0);
     Control              : std_logic_vector(31 downto 0);
     IrqFlag              : std_logic_vector(31 downto 0);
     IrqEnable            : std_logic_vector(31 downto 0);
     PulseIrqMap          : std_logic_vector(31 downto 0);
     SWEvent              : std_logic_vector(31 downto 0);
     DataBufCtrl          : std_logic_vector(31 downto 0);
     TXDataBufCtrl        : std_logic_vector(31 downto 0);
     TxSegBufCtrl         : std_logic_vector(31 downto 0);
     FWVersion            : std_logic_vector(31 downto 0);
     EvCntPresc           : std_logic_vector(31 downto 0);
     UsecDivider          : std_logic_vector(31 downto 0);
     ClockControl         : std_logic_vector(31 downto 0);
     SecSR                : std_logic_vector(31 downto 0);
     SecCounter           : std_logic_vector(31 downto 0);
     EventCounter         : std_logic_vector(31 downto 0);
     SecLatch             : std_logic_vector(31 downto 0);
     EvCntLatch           : std_logic_vector(31 downto 0);
     EvFIFOSec            : std_logic_vector(31 downto 0);
     EvFIFOEvCnt          : std_logic_vector(31 downto 0);
     EvFIFOCode           : std_logic_vector(31 downto 0);
     LogStatus            : std_logic_vector(31 downto 0);
     GPIODir              : std_logic_vector(31 downto 0);
     GPIOIn               : std_logic_vector(31 downto 0);
     GPIOOut              : std_logic_vector(31 downto 0);
     DCTarget             : std_logic_vector(31 downto 0);
     DCRxValue            : std_logic_vector(31 downto 0);
     DCIntValue           : std_logic_vector(31 downto 0);
     DCStatus             : std_logic_vector(31 downto 0);
     TopologyID           : std_logic_vector(31 downto 0);
     SeqRamCtrl           : std_logic_vector(31 downto 0);
     Prescaler0           : std_logic_vector(31 downto 0);
     Prescaler1           : std_logic_vector(31 downto 0);
     Prescaler2           : std_logic_vector(31 downto 0);
     Prescaler3           : std_logic_vector(31 downto 0);
     Prescaler4           : std_logic_vector(31 downto 0);
     Prescaler5           : std_logic_vector(31 downto 0);
     Prescaler6           : std_logic_vector(31 downto 0);
     Prescaler7           : std_logic_vector(31 downto 0);
     PrescPhase0          : std_logic_vector(31 downto 0);
     PrescPhase1          : std_logic_vector(31 downto 0);
     PrescPhase2          : std_logic_vector(31 downto 0);
     PrescPhase3          : std_logic_vector(31 downto 0);
     PrescPhase4          : std_logic_vector(31 downto 0);
     PrescPhase5          : std_logic_vector(31 downto 0);
     PrescPhase6          : std_logic_vector(31 downto 0);
     PrescPhase7          : std_logic_vector(31 downto 0);
     PrescTrig0           : std_logic_vector(31 downto 0);
     PrescTrig1           : std_logic_vector(31 downto 0);
     PrescTrig2           : std_logic_vector(31 downto 0);
     PrescTrig3           : std_logic_vector(31 downto 0);
     PrescTrig4           : std_logic_vector(31 downto 0);
     PrescTrig5           : std_logic_vector(31 downto 0);
     PrescTrig6           : std_logic_vector(31 downto 0);
     PrescTrig7           : std_logic_vector(31 downto 0);
     DBusTrig0            : std_logic_vector(31 downto 0);
     DBusTrig1            : std_logic_vector(31 downto 0);
     DBusTrig2            : std_logic_vector(31 downto 0);
     DBusTrig3            : std_logic_vector(31 downto 0);
     DBusTrig4            : std_logic_vector(31 downto 0);
     DBusTrig5            : std_logic_vector(31 downto 0);
     DBusTrig6            : std_logic_vector(31 downto 0);
     DBusTrig7            : std_logic_vector(31 downto 0);
     Pulse0Ctrl           : std_logic_vector(31 downto 0);
     Pulse0Presc          : std_logic_vector(31 downto 0);
     Pulse0Delay          : std_logic_vector(31 downto 0);
     Pulse0Width          : std_logic_vector(31 downto 0);
     Pulse1Ctrl           : std_logic_vector(31 downto 0);
     Pulse1Presc          : std_logic_vector(31 downto 0);
     Pulse1Delay          : std_logic_vector(31 downto 0);
     Pulse1Width          : std_logic_vector(31 downto 0);
     Pulse2Ctrl           : std_logic_vector(31 downto 0);
     Pulse2Presc          : std_logic_vector(31 downto 0);
     Pulse2Delay          : std_logic_vector(31 downto 0);
     Pulse2Width          : std_logic_vector(31 downto 0);
     Pulse3Ctrl           : std_logic_vector(31 downto 0);
     Pulse3Presc          : std_logic_vector(31 downto 0);
     Pulse3Delay          : std_logic_vector(31 downto 0);
     Pulse3Width          : std_logic_vector(31 downto 0);
     Pulse4Ctrl           : std_logic_vector(31 downto 0);
     Pulse4Presc          : std_logic_vector(31 downto 0);
     Pulse4Delay          : std_logic_vector(31 downto 0);
     Pulse4Width          : std_logic_vector(31 downto 0);
     Pulse5Ctrl           : std_logic_vector(31 downto 0);
     Pulse5Presc          : std_logic_vector(31 downto 0);
     Pulse5Delay          : std_logic_vector(31 downto 0);
     Pulse5Width          : std_logic_vector(31 downto 0);
     Pulse6Ctrl           : std_logic_vector(31 downto 0);
     Pulse6Presc          : std_logic_vector(31 downto 0);
     Pulse6Delay          : std_logic_vector(31 downto 0);
     Pulse6Width          : std_logic_vector(31 downto 0);
     Pulse7Ctrl           : std_logic_vector(31 downto 0);
     Pulse7Presc          : std_logic_vector(31 downto 0);
     Pulse7Delay          : std_logic_vector(31 downto 0);
     Pulse7Width          : std_logic_vector(31 downto 0);
     Pulse8Ctrl           : std_logic_vector(31 downto 0);
     Pulse8Presc          : std_logic_vector(31 downto 0);
     Pulse8Delay          : std_logic_vector(31 downto 0);
     Pulse8Width          : std_logic_vector(31 downto 0);
     Pulse9Ctrl           : std_logic_vector(31 downto 0);
     Pulse9Presc          : std_logic_vector(31 downto 0);
     Pulse9Delay          : std_logic_vector(31 downto 0);
     Pulse9Width          : std_logic_vector(31 downto 0);
     Pulse10Ctrl          : std_logic_vector(31 downto 0);
     Pulse10Presc         : std_logic_vector(31 downto 0);
     Pulse10Delay         : std_logic_vector(31 downto 0);
     Pulse10Width         : std_logic_vector(31 downto 0);
     Pulse11Ctrl          : std_logic_vector(31 downto 0);
     Pulse11Presc         : std_logic_vector(31 downto 0);
     Pulse11Delay         : std_logic_vector(31 downto 0);
     Pulse11Width         : std_logic_vector(31 downto 0);
     Pulse12Ctrl          : std_logic_vector(31 downto 0);
     Pulse12Presc         : std_logic_vector(31 downto 0);
     Pulse12Delay         : std_logic_vector(31 downto 0);
     Pulse12Width         : std_logic_vector(31 downto 0);
     Pulse13Ctrl          : std_logic_vector(31 downto 0);
     Pulse13Presc         : std_logic_vector(31 downto 0);
     Pulse13Delay         : std_logic_vector(31 downto 0);
     Pulse13Width         : std_logic_vector(31 downto 0);
     Pulse14Ctrl          : std_logic_vector(31 downto 0);
     Pulse14Presc         : std_logic_vector(31 downto 0);
     Pulse14Delay         : std_logic_vector(31 downto 0);
     Pulse14Width         : std_logic_vector(31 downto 0);
     Pulse15Ctrl          : std_logic_vector(31 downto 0);
     Pulse15Presc         : std_logic_vector(31 downto 0);
     Pulse15Delay         : std_logic_vector(31 downto 0);
     Pulse15Width         : std_logic_vector(31 downto 0);
     Pulse16Ctrl          : std_logic_vector(31 downto 0);
     Pulse16Presc         : std_logic_vector(31 downto 0);
     Pulse16Delay         : std_logic_vector(31 downto 0);
     Pulse16Width         : std_logic_vector(31 downto 0);
     Pulse17Ctrl          : std_logic_vector(31 downto 0);
     Pulse17Presc         : std_logic_vector(31 downto 0);
     Pulse17Delay         : std_logic_vector(31 downto 0);
     Pulse17Width         : std_logic_vector(31 downto 0);
     Pulse18Ctrl          : std_logic_vector(31 downto 0);
     Pulse18Presc         : std_logic_vector(31 downto 0);
     Pulse18Delay         : std_logic_vector(31 downto 0);
     Pulse18Width         : std_logic_vector(31 downto 0);
     Pulse19Ctrl          : std_logic_vector(31 downto 0);
     Pulse19Presc         : std_logic_vector(31 downto 0);
     Pulse19Delay         : std_logic_vector(31 downto 0);
     Pulse19Width         : std_logic_vector(31 downto 0);
     Pulse20Ctrl          : std_logic_vector(31 downto 0);
     Pulse20Presc         : std_logic_vector(31 downto 0);
     Pulse20Delay         : std_logic_vector(31 downto 0);
     Pulse20Width         : std_logic_vector(31 downto 0);
     Pulse21Ctrl          : std_logic_vector(31 downto 0);
     Pulse21Presc         : std_logic_vector(31 downto 0);
     Pulse21Delay         : std_logic_vector(31 downto 0);
     Pulse21Width         : std_logic_vector(31 downto 0);
     Pulse22Ctrl          : std_logic_vector(31 downto 0);
     Pulse22Presc         : std_logic_vector(31 downto 0);
     Pulse22Delay         : std_logic_vector(31 downto 0);
     Pulse22Width         : std_logic_vector(31 downto 0);
     Pulse23Ctrl          : std_logic_vector(31 downto 0);
     Pulse23Presc         : std_logic_vector(31 downto 0);
     Pulse23Delay         : std_logic_vector(31 downto 0);
     Pulse23Width         : std_logic_vector(31 downto 0);
     Pulse24Ctrl          : std_logic_vector(31 downto 0);
     Pulse24Presc         : std_logic_vector(31 downto 0);
     Pulse24Delay         : std_logic_vector(31 downto 0);
     Pulse24Width         : std_logic_vector(31 downto 0);
     Pulse25Ctrl          : std_logic_vector(31 downto 0);
     Pulse25Presc         : std_logic_vector(31 downto 0);
     Pulse25Delay         : std_logic_vector(31 downto 0);
     Pulse25Width         : std_logic_vector(31 downto 0);
     Pulse26Ctrl          : std_logic_vector(31 downto 0);
     Pulse26Presc         : std_logic_vector(31 downto 0);
     Pulse26Delay         : std_logic_vector(31 downto 0);
     Pulse26Width         : std_logic_vector(31 downto 0);
     Pulse27Ctrl          : std_logic_vector(31 downto 0);
     Pulse27Presc         : std_logic_vector(31 downto 0);
     Pulse27Delay         : std_logic_vector(31 downto 0);
     Pulse27Width         : std_logic_vector(31 downto 0);
     Pulse28Ctrl          : std_logic_vector(31 downto 0);
     Pulse28Presc         : std_logic_vector(31 downto 0);
     Pulse28Delay         : std_logic_vector(31 downto 0);
     Pulse28Width         : std_logic_vector(31 downto 0);
     Pulse29Ctrl          : std_logic_vector(31 downto 0);
     Pulse29Presc         : std_logic_vector(31 downto 0);
     Pulse29Delay         : std_logic_vector(31 downto 0);
     Pulse29Width         : std_logic_vector(31 downto 0);
     Pulse30Ctrl          : std_logic_vector(31 downto 0);
     Pulse30Presc         : std_logic_vector(31 downto 0);
     Pulse30Delay         : std_logic_vector(31 downto 0);
     Pulse30Width         : std_logic_vector(31 downto 0);
     Pulse31Ctrl          : std_logic_vector(31 downto 0);
     Pulse31Presc         : std_logic_vector(31 downto 0);
     Pulse31Delay         : std_logic_vector(31 downto 0);
     Pulse31Width         : std_logic_vector(31 downto 0);
     ESSStatus            : std_logic_vector(31 downto 0);
     ESSControl           : std_logic_vector(31 downto 0);
     ESSExtSecCounter     : std_logic_vector(31 downto 0);
     ESSExtEventCounter   : std_logic_vector(31 downto 0);
  end record;

  type transfer_shadow_group_t is record
    none : std_logic;
  end record;


  

end register_bank_config;
